package fsm_pkg is
    type fsm_state is
    (
        START,
        S0,
        S1,
        S2
    );
end package fsm_pkg;